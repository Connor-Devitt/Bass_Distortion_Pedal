** Profile: "SCHEMATIC1-Freq_Sweep"  [ e:\user\connor\documents\ee projects\distortion_pedal\bass_distortion_pedal\electrical\simulation\distortion_pedal_sim-PSpiceFiles\SCHEMATIC1\Freq_Sweep.sim ] 

** Creating circuit file "Freq_Sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Connor\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 1000 40Hz 20KHz
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
