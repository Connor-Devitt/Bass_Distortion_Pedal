** Profile: "SCHEMATIC1-balance_sweep"  [ e:\user\connor\documents\ee projects\distortion_pedal\bass_distortion_pedal\electrical\simulation\distortion_pedal_sim-PSpiceFiles\SCHEMATIC1\balance_sweep.sim ] 

** Creating circuit file "balance_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Connor\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 50ms 0 0.001ms 
.STEP LIN PARAM set_pot3 5k 45k 5k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
